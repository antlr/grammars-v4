module top;
  initial $system("mv design.v adder.v");
endmodule
