../../vhdl/examples/standard.vhd