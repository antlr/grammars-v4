task automatic show(const ref byte data[]);
  for (int j = 0; j < data.size; j++) $display(data[j]);
endtask
