../../vhdl/examples/numeric_std.vhd