../../vhdl/examples/unsigned.vhd