typedef struct {
  int addr = 1 + constant;
  int crc;
  byte data[4] = '{4{1}};
} packet1;
