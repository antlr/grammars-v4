../../vhdl/examples/textio.vhd