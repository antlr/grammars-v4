module test;
  logic clk;
  logic a, b;
  logic c, d;
endmodule
