../../vhdl/examples/signed.vhd