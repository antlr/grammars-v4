task t;
  logic s;
  begin : b
    logic r;
    t.b.r = 0;
    b.r = 0;
    r = 0;
    t.s = 0;
    s = 0;
  end
endtask
