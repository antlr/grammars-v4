../../vhdl/examples/std_logic_1164.vhd