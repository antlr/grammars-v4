module m (
    input clock
);
  logic a;
endmodule : m
