struct {
  bit [7:0] A;
  bit [7:0] B;
  byte C;
} abc;
