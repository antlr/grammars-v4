../../vhdl/examples/std_logic_1164_body.vhd