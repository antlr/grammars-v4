../../vhdl/examples/numeric_std-body.vhd