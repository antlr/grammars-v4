../../vhdl/examples/std_logic_textio.vhd