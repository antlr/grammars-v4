class C #(
    int p = 1
);
  parameter int q = 5;
  static task t;
    int p;
    int x = C::p;
  endtask
endclass
