../../vhdl/examples/misc.vhd