module top (a);
  input a;
  wire hello;
  NOT u1 (hello, a);
endmodule
