module m;
  import q::*;
  wire a = c;
  import p::c;
endmodule
