../../vhdl/examples/add_pkg.vhd