../../vhdl/examples/arith.vhd