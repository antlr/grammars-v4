../../vhdl/examples/numeric_bit-body.vhd