module test (
    input [7:0] a,
    input signed [7:0] b,
    c,
    d,
    output [7:0] e,
    output var signed [7:0] f,
    g,
    output signed [7:0] h
);
endmodule
module cpuMod (
    interface d,
    interface j
);
endmodule
