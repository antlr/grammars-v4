task task1(integer a, obj_example myexample);
  if (myexample == null) myexample = new;
endtask
