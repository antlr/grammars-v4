../../vhdl/examples/numeric_bit.vhd